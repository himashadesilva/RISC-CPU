module datapath(input_addr,instruction);
input [3:0] input_addr;
output reg [31:0] instruction;

wire[3:0] current_addr;
wire [



endmodule
